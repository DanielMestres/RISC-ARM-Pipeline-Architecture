module IDEX_Register (
    
);