module Adder (

);