// This module is to initialize and connect everything
// Create clk here
// Takes no input nor produces any outputs

module main;