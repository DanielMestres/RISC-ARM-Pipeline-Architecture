module MEMWB_Register (
    
);