module Condition_Handler (

);