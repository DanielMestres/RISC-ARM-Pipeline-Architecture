module EXMEM_Register (
    output reg size_o,
    output reg enable_o,
    output reg rw_o,
    output reg  load_o,
    output reg rf_o,
    input size_i,
    input enable_i,
    input rw_i,
    input load_i,
    input rf_i,
    input CLK,
    input CLR
);

    always@(posedge CLK) begin
        if(CLR) begin
        load_o = 1'b0;
        rf_o = 1'b0;
        size_o = 1'b0;
        enable_o = 1'b0;
        rw_o = 1'b0;
        end else begin
            load_o = load_i;
            rf_o = rf_i;
            size_o = size_i;
            enable_o = enable_i;
            rw_o = rw_i;
        end
    end
endmodule