module PC_4_Adder (

);