module EXMEM_Register (
    
);