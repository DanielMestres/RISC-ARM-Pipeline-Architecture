module Mux (

);