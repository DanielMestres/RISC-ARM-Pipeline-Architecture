module Mux_4_1 (

);