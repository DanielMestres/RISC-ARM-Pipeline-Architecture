module IFID_Register (
    
);