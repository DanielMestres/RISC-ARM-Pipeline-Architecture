module RAM (
  
  );

  always @(*) begin
    
  end
endmodule