module Hazard_Unit (

);