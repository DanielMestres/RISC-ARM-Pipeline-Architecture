module Control_Unit (
    input [31:0] IR_in,
    output SE_ID_out,
    output LI_ID_out,
    output RF_ID_out,
    output B_ID_out,
    output [3:0] opcode_out
);
endmodule